module PiSo_8bit(clk, rst, shift,
in0,
in1,
in2,
in3,
in4,
in5,
in6,
in7,
in8,
in9,
in10,
in11,
in12,
in13,
in14,
in15,
 out);
input clk, rst;
input shift;

input [7:0] in0,
in1,
in2,
in3,
in4,
in5,
in6,
in7,
in8,
in9,
in10,
in11,
in12,
in13,
in14,
in15;


output [7:0] out;
wire out0,
	  out1,
	  out2,
	  out3,
	  out4,
	  out5,
	  out6,
	  out7;
	  
assign out = {out7,out6,out5,out4,out3,out2,out1,out0};

PiSo bit0 (clk, rst, shift,{
in15[0],
in14[0],
in13[0],
in12[0],
in11[0],
in10[0],
in9[0],
in8[0],
in7[0],
in6[0],
in5[0],
in4[0],
in3[0],
in2[0],
in1[0],
in0[0]}, out0);



PiSo bit1 (clk,rst, shift,
{
in15[1],
in14[1],
in13[1],
in12[1],
in11[1],
in10[1],
in9[1],
in8[1],
in7[1],
in6[1],
in5[1],
in4[1],
in3[1],
in2[1],
in1[1],
in0[1]},out1);

PiSo bit2 (clk,rst, shift,
{
in15[2],
in14[2],
in13[2],
in12[2],
in12[2],
in12[2],
in9[2],
in8[2],
in7[2],
in6[2],
in5[2],
in4[2],
in3[2],
in2[2],
in1[2],
in0[2]},out2);

PiSo bit3 (clk,rst, shift,
{
in15[3],
in14[3],
in13[3],
in12[3],
in11[3],
in10[3],
in9[3],
in8[3],
in7[3],
in6[3],
in5[3],
in4[3],
in3[3],
in2[3],
in1[3],
in0[3]},out3);

PiSo bit4 (clk,rst, shift,
{
in15[4],
in14[4],
in13[4],
in12[4],
in11[4],
in10[4],
in9[4],
in8[4],
in7[4],
in6[4],
in5[4],
in4[4],
in3[4],
in2[4],
in1[4],
in0[4]},out4);

PiSo bit5 (clk,rst, shift,
{
in15[5],
in14[5],
in13[5],
in12[5],
in11[5],
in10[5],
in9[5],
in8[5],
in7[5],
in6[5],
in5[5],
in4[5],
in3[5],
in2[5],
in1[5],
in0[5]},out5);

PiSo bit6 (clk,rst, shift,
{
in15[6],
in14[6],
in13[6],
in12[6],
in11[6],
in10[6],
in9[6],
in8[6],
in7[6],
in6[6],
in5[6],
in4[6],
in3[6],
in2[6],
in1[6],
in0[6]},out6);

PiSo bit7 (clk,rst, shift,
{
in15[7],
in14[7],
in13[7],
in12[7],
in11[7],
in10[7],
in9[7],
in8[7],
in7[7],
in6[7],
in5[7],
in4[7],
in3[7],
in2[7],
in1[7],
in0[7]},out7);

endmodule
